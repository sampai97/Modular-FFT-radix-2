library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package twiddle_type_pkg is
constant N_bit : integer := 15;         --sample depth
constant N_twiddle : integer := 192;    --number of twiddle factor, need to change if change number of points
type twiddle_vector is array (0 to N_twiddle-1) of signed(N_bit-1 downto 0);

constant twiddle_re : twiddle_vector := ("010000000000000", --real part
"001111111011001",
"001111101100011",
"001111010011111",
"001110110010000",
"001110000111001",
"001101010011011",
"001100010111101",
"001011010100001",
"001010001001101",
"001000111000111",
"000111100010110",
"000110000111111",
"000100101001010",
"000011000111110",
"000001100100011",
"000000000000000",
"111110011011101",
"111100111000010",
"111011010110110",
"111001111000001",
"111000011101010",
"110111000111001",
"110101110110011",
"110100101011111",
"110011101000011",
"110010101100101",
"110001111000111",
"110001001110000",
"110000101100001",
"110000010011101",
"110000000100111",
"010000000000000",
"001111101100011",
"001110110010000",
"001101010011011",
"001011010100001",
"001000111000111",
"000110000111111",
"000011000111110",
"000000000000000",
"111100111000010",
"111001111000001",
"110111000111001",
"110100101011111",
"110010101100101",
"110001001110000",
"110000010011101",
"010000000000000",
"001111101100011",
"001110110010000",
"001101010011011",
"001011010100001",
"001000111000111",
"000110000111111",
"000011000111110",
"000000000000000",
"111100111000010",
"111001111000001",
"110111000111001",
"110100101011111",
"110010101100101",
"110001001110000",
"110000010011101",
"010000000000000",
"001110110010000",
"001011010100001",
"000110000111111",
"000000000000000",
"111001111000001",
"110100101011111",
"110001001110000",
"010000000000000",
"001110110010000",
"001011010100001",
"000110000111111",
"000000000000000",
"111001111000001",
"110100101011111",
"110001001110000",
"010000000000000",
"001110110010000",
"001011010100001",
"000110000111111",
"000000000000000",
"111001111000001",
"110100101011111",
"110001001110000",
"010000000000000",
"001110110010000",
"001011010100001",
"000110000111111",
"000000000000000",
"111001111000001",
"110100101011111",
"110001001110000",
"010000000000000",
"001011010100001",
"000000000000000",
"110100101011111",
"010000000000000",
"001011010100001",
"000000000000000",
"110100101011111",
"010000000000000",
"001011010100001",
"000000000000000",
"110100101011111",
"010000000000000",
"001011010100001",
"000000000000000",
"110100101011111",
"010000000000000",
"001011010100001",
"000000000000000",
"110100101011111",
"010000000000000",
"001011010100001",
"000000000000000",
"110100101011111",
"010000000000000",
"001011010100001",
"000000000000000",
"110100101011111",
"010000000000000",
"001011010100001",
"000000000000000",
"110100101011111",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"000000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000",
"010000000000000");

constant twiddle_im : twiddle_vector := ("000000000000000", --imagginary part
"111110011011101",
"111100111000010",
"111011010110110",
"111001111000001",
"111000011101010",
"110111000111001",
"110101110110011",
"110100101011111",
"110011101000011",
"110010101100101",
"110001111000111",
"110001001110000",
"110000101100001",
"110000010011101",
"110000000100111",
"110000000000000",
"110000000100111",
"110000010011101",
"110000101100001",
"110001001110000",
"110001111000111",
"110010101100101",
"110011101000011",
"110100101011111",
"110101110110011",
"110111000111001",
"111000011101010",
"111001111000001",
"111011010110110",
"111100111000010",
"111110011011101",
"000000000000000",
"111100111000010",
"111001111000001",
"110111000111001",
"110100101011111",
"110010101100101",
"110001001110000",
"110000010011101",
"110000000000000",
"110000010011101",
"110001001110000",
"110010101100101",
"110100101011111",
"110111000111001",
"111001111000001",
"111100111000010",
"000000000000000",
"111100111000010",
"111001111000001",
"110111000111001",
"110100101011111",
"110010101100101",
"110001001110000",
"110000010011101",
"110000000000000",
"110000010011101",
"110001001110000",
"110010101100101",
"110100101011111",
"110111000111001",
"111001111000001",
"111100111000010",
"000000000000000",
"111001111000001",
"110100101011111",
"110001001110000",
"110000000000000",
"110001001110000",
"110100101011111",
"111001111000001",
"000000000000000",
"111001111000001",
"110100101011111",
"110001001110000",
"110000000000000",
"110001001110000",
"110100101011111",
"111001111000001",
"000000000000000",
"111001111000001",
"110100101011111",
"110001001110000",
"110000000000000",
"110001001110000",
"110100101011111",
"111001111000001",
"000000000000000",
"111001111000001",
"110100101011111",
"110001001110000",
"110000000000000",
"110001001110000",
"110100101011111",
"111001111000001",
"000000000000000",
"110100101011111",
"110000000000000",
"110100101011111",
"000000000000000",
"110100101011111",
"110000000000000",
"110100101011111",
"000000000000000",
"110100101011111",
"110000000000000",
"110100101011111",
"000000000000000",
"110100101011111",
"110000000000000",
"110100101011111",
"000000000000000",
"110100101011111",
"110000000000000",
"110100101011111",
"000000000000000",
"110100101011111",
"110000000000000",
"110100101011111",
"000000000000000",
"110100101011111",
"110000000000000",
"110100101011111",
"000000000000000",
"110100101011111",
"110000000000000",
"110100101011111",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"110000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000",
"000000000000000");
end package twiddle_type_pkg;
